`undef BITWIDTH
