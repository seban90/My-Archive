`define BITWIDTH 8
