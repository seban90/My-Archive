`timescale 1ns/1ps

module t;
	`include "clock_reset.vinc"
	`include "pkg.vinc"
endmodule
