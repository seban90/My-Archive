`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module half_adder_structural(din1, din2, sum, carry);

    input din1, din2;
    output sum, carry;
     
    xor (sum, din1, din2);
    and (carry, din1, din2);
     
endmodule
